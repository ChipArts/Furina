// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : InstructionFetchUnit.sv
// Create  : 2024-03-01 16:11:09
// Revise  : 2024-03-01 16:11:09
// Description :
//   取指单元
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ...
// ==============================================================================

`include "InstructionFetchUnit.svh"

module InstructionFetchUnit (
  input clk,    // Clock
  input a_rst_n,  // Asynchronous reset active low
  
);

endmodule : InstructionFetchUnit


