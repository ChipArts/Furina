// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : CSR.svh
// Create  : 2024-03-18 22:28:51
// Revise  : 2024-03-18 22:31:58
// Description :
//   ...
//   ...
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ...
// ==============================================================================

`ifndef _CSR_SVH_
`define _CSR_SVH_

typedef logic[5:0] ExceptionType;

`define EXC_NONE (6'd0)



`endif  // _CSR_SVH_