// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : AXI4.sv
// Create  : 2024-01-13 20:29:55
// Revise  : 2024-01-13 20:29:55
// Description :
//    An AXI4(Advanced eXtensible Interface) interface.
// Parameter   :
//    ...
//    ...
// IO Port     :
//    ...
//    ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// 24-01-13 |            |     0.1     |    Original Version
// ==============================================================================

interface AXI4 #(
  parameter int unsigned AXI_ADDR_WIDTH  = 32,
  parameter int unsigned AXI_DATA_WIDTH  = 32,
  parameter int unsigned AXI_ID_WIDTH    = 4,
  parameter int unsigned AXI_USER_WIDTH  = 1
);

  localparam int unsigned AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
  
  typedef logic [AXI_ID_WIDTH-1:0]   id_t;
  typedef logic [AXI_ADDR_WIDTH-1:0] addr_t;
  typedef logic [AXI_DATA_WIDTH-1:0] data_t;
  typedef logic [AXI_STRB_WIDTH-1:0] strb_t;
  typedef logic [AXI_USER_WIDTH-1:0] user_t;
  typedef logic [4             -1:0] len_t;
  typedef logic [3             -1:0] size_t;
  typedef logic [2             -1:0] burst_t;
  typedef logic [4             -1:0] cache_t;
  typedef logic [3             -1:0] prot_t;
  typedef logic [1             -1:0] qos_t;
  typedef logic [1             -1:0] region_t;
  typedef logic [1             -1:0] resp_t;
  
  id_t     aw_id;
  addr_t   aw_addr;
  len_t    aw_len;
  size_t   aw_size;
  burst_t  aw_burst;
  logic    aw_lock;
  cache_t  aw_cache;
  prot_t   aw_prot;
  qos_t    aw_qos;
  region_t aw_region;
  user_t   aw_user;
  logic    aw_valid;
  logic    aw_ready;
  
  id_t     w_id;
  data_t   w_data;
  strb_t   w_strb;
  logic    w_last;
  user_t   w_user;
  logic    w_valid;
  logic    w_ready;
  
  id_t     b_id;
  resp_t   b_resp;
  user_t   b_user;
  logic    b_valid;
  logic    b_ready;
  
  id_t     ar_id;
  addr_t   ar_addr;
  len_t    ar_len;
  size_t   ar_size;
  burst_t  ar_burst;
  logic    ar_lock;
  cache_t  ar_cache;
  prot_t   ar_prot;
  qos_t    ar_qos;
  region_t ar_region;
  user_t   ar_user;
  logic    ar_valid;
  logic    ar_ready;
  
  id_t     r_id;
  data_t   r_data;
  resp_t   r_resp;
  logic    r_last;
  user_t   r_user;
  logic    r_valid;
  logic    r_ready;
  
  modport Master (
    output aw_id, aw_addr, aw_len, aw_size, aw_burst, aw_lock, aw_cache, aw_prot, aw_qos, aw_region, aw_user, aw_valid, input aw_ready,
    output w_id, w_data, w_strb, w_last, w_user, w_valid, input w_ready,
    input b_id, b_resp, b_user, b_valid, output b_ready,
    output ar_id, ar_addr, ar_len, ar_size, ar_burst, ar_lock, ar_cache, ar_prot, ar_qos, ar_region, ar_user, ar_valid, input ar_ready,
    input r_id, r_data, r_resp, r_last, r_user, r_valid, output r_ready
  );
  
  modport Slave (
    input aw_id, aw_addr, aw_len, aw_size, aw_burst, aw_lock, aw_cache, aw_prot, aw_qos, aw_region, aw_user, aw_valid, output aw_ready,
    input w_id, w_data, w_strb, w_last, w_user, w_valid, output w_ready,
    output b_id, b_resp, b_user, b_valid, input b_ready,
    input ar_id, ar_addr, ar_len, ar_size, ar_burst, ar_lock, ar_cache, ar_prot, ar_qos, ar_region, ar_user, ar_valid, output ar_ready,
    output r_id, r_data, r_resp, r_last, r_user, r_valid, input r_ready
  );
  
  modport Monitor (
    input aw_id, aw_addr, aw_len, aw_size, aw_burst, aw_lock, aw_cache, aw_prot, aw_qos, aw_region, aw_user, aw_valid, aw_ready,
        w_id, w_data, w_strb, w_last, w_user, w_valid, w_ready,
        b_id, b_resp, b_user, b_valid, b_ready,
        ar_id, ar_addr, ar_len, ar_size, ar_burst, ar_lock, ar_cache, ar_prot, ar_qos, ar_region, ar_user, ar_valid, ar_ready,
        r_id, r_data, r_resp, r_last, r_user, r_valid, r_ready
  );

endinterface
