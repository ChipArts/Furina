// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : FetchAddressQueue.sv
// Create  : 2024-02-12 16:37:58
// Revise  : 2024-02-13 11:32:13
// Description :
//   ...
//   ...
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ...
// ==============================================================================

`include "config.svh"
`include "common.svh"
`include "bpu.svh"

module FetchAddressQueue (
  input clk,    // Clock
  input rst_n,  // Asynchronous reset active low
  input BPU2FAQSt bpu2faq_st_i,
);

endmodule : FetchAddressQueue