// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : MemoryBlock.sv
// Create  : 2024-03-17 22:34:12
// Revise  : 2024-03-20 23:17:26
// Description :
//   ...
//   ...
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ...
// ==============================================================================

`include "config.svh"
`include "Decoder.svh"

module MemoryBlock (
  input clk,    // Clock
  input rst_n,  // Asynchronous reset active low
  
);

endmodule : MemoryBlock

