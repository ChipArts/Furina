// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : Decoder.sv
// Create  : 2024-03-01 16:02:44
// Revise  : 2024-03-01 16:02:44
// Description :
//   解码器
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ==============================================================================

`include "Decoder.svh"

module Decoder (
  input logic [31:0] instr,
  output OptionCodeSt option_code
);

  // TODO: generate decoder by SpinalHDL

endmodule : Decoder
