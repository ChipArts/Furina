// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : MemoryBlock.sv
// Create  : 2024-03-17 22:34:12
// Revise  : 2024-03-27 20:36:24
// Description :
//   ...
//   ...
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ...
// ==============================================================================

`include "config.svh"
`include "common.svh"
`include "Decoder.svh"
`include "Pipeline.svh"
`include "MemoryManagementUnit.svh"

module MemoryBlock (
  input clk,    // Clock
  input a_rst_n,  // Asynchronous reset active low
  input flush_i,
  /* exe */
  input MemExeSt exe_i,
  output logic exe_ready_o,
  /* other exe io */
  output MmuAddrTransReqSt addr_trans_req,
  input MmuAddrTransRspSt addr_trans_rsp,
  AXI4.Master axi4_mst,
  /* wirte back */
  output MemWbSt wb_o,
  input logic wb_ready_i
);

  `RESET_LOGIC(clk, a_rst_n, rst_n);
  logic s0_ready, s1_ready;

/*================================== stage0 ===================================*/
  // regfile comb输出 数据缓存一拍
  always_comb begin
    s0_ready = s1_ready;
  end


/*================================== stage1 ===================================*/
  // TODO: exe cacop micro
  MemExeSt s1_exe;

  always_ff @(posedge clk or negedge rst_n) begin
    if(~rst_n || flush_i) begin
      s1_exe <= '0;
    end else begin
      if (s1_ready) begin
        s1_exe <= exe_i;
      end
    end
  end

  DCacheReqSt dcache_req;
  DCacheRspSt dcache_rsp;
  MmuAddrTransReqSt dcache_addr_trans_req;
  MmuAddrTransRspSt dcache_addr_trans_rsp;

  always_comb begin
    s1_ready = dcache_rsp.ready | ~s1_exe.base.valid;

    dcache_req.valid = s1_exe.base.valid;
    dcache_req.ready = '1;
    dcache_req.vaddr = s1_exe.base.src0 + s1_exe.imm;
    dcache_req.wdata = s1_exe.base.src1;
    dcache_req.rob_idx = s1_exe.base.rob_idx;
    dcache_req.align_op = s1_exe.mem_oc.align_op;
    dcache_req.mem_type = s1_exe.mem_oc.mem_type;

    
    addr_trans_req = dcache_addr_trans_req;
    dcache_addr_trans_rsp = addr_trans_rsp;
  end

  // DCache视为一个多周期的模块
  DCache inst_DCache
  (
    .clk              (clk),
    .a_rst_n          (rst_n),
    .flush_i          (flush_i),
    .req              (dcache_req),
    .rsp              (dcache_rsp),
    .addr_trans_req   (dcache_addr_trans_req),
    .addr_trans_rsp   (dcache_addr_trans_rsp),
    .axi4_mst         (axi4_mst)
  );

/*================================== stage2 ===================================*/
  // 产生commit信息
  always_comb begin
    wb_o.base.valid = dcache_rsp.valid;
    wb_o.base.we = dcache_rsp.mem_type == `MEM_LOAD;
    wb_o.base.wdata = dcache_rsp.rdata;
    wb_o.base.rob_idx = dcache_rsp.rob_idx;
    wb_o.base.pdest = dcache_rsp.pdest;
    wb_o.base.exception = dcache_rsp.exception;
    wb_o.base.ecode = dcache_rsp.ecode;
  end


endmodule : MemoryBlock

