// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : Decoder.sv
// Create  : 2024-03-01 16:02:44
// Revise  : 2024-03-01 16:02:44
// Description :
//   解码器
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ==============================================================================

`include "Decoder.svh"

// Generator : SpinalHDL v1.10.1    git head : 2527c7c6b0fb0f95e5e1a5722a0be732b364ce43
// Component : Decoder
// Git hash  : d174bcf88ffe8bc86a1212f21a64337548cbeb1c

`timescale 1ns/1ps

module Decoder (
  input  wire [31:0]   instr_i,
  output wire [58:0]   option_code_o
);

  wire       [31:0]   _zz_ctrl;
  wire                _zz_ctrl_1;
  wire       [0:0]    _zz_ctrl_2;
  wire       [31:0]   _zz_ctrl_3;
  wire       [3:0]    _zz_ctrl_4;
  wire       [31:0]   _zz_ctrl_5;
  wire       [31:0]   _zz_ctrl_6;
  wire                _zz_ctrl_7;
  wire       [31:0]   _zz_ctrl_8;
  wire       [0:0]    _zz_ctrl_9;
  wire       [31:0]   _zz_ctrl_10;
  wire       [31:0]   _zz_ctrl_11;
  wire       [0:0]    _zz_ctrl_12;
  wire       [31:0]   _zz_ctrl_13;
  wire       [31:0]   _zz_ctrl_14;
  wire       [0:0]    _zz_ctrl_15;
  wire       [31:0]   _zz_ctrl_16;
  wire       [0:0]    _zz_ctrl_17;
  wire       [31:0]   _zz_ctrl_18;
  wire       [0:0]    _zz_ctrl_19;
  wire       [31:0]   _zz_ctrl_20;
  wire                _zz_ctrl_21;
  wire                _zz_ctrl_22;
  wire       [31:0]   _zz_ctrl_23;
  wire                _zz_ctrl_24;
  wire       [31:0]   _zz_ctrl_25;
  wire       [0:0]    _zz_ctrl_26;
  wire                _zz_ctrl_27;
  wire       [31:0]   _zz_ctrl_28;
  wire       [19:0]   _zz_ctrl_29;
  wire       [2:0]    _zz_ctrl_30;
  wire                _zz_ctrl_31;
  wire       [31:0]   _zz_ctrl_32;
  wire       [0:0]    _zz_ctrl_33;
  wire       [31:0]   _zz_ctrl_34;
  wire       [31:0]   _zz_ctrl_35;
  wire       [0:0]    _zz_ctrl_36;
  wire       [31:0]   _zz_ctrl_37;
  wire       [31:0]   _zz_ctrl_38;
  wire                _zz_ctrl_39;
  wire       [0:0]    _zz_ctrl_40;
  wire       [31:0]   _zz_ctrl_41;
  wire       [31:0]   _zz_ctrl_42;
  wire       [2:0]    _zz_ctrl_43;
  wire                _zz_ctrl_44;
  wire       [31:0]   _zz_ctrl_45;
  wire       [0:0]    _zz_ctrl_46;
  wire       [31:0]   _zz_ctrl_47;
  wire       [31:0]   _zz_ctrl_48;
  wire       [0:0]    _zz_ctrl_49;
  wire       [31:0]   _zz_ctrl_50;
  wire       [31:0]   _zz_ctrl_51;
  wire       [0:0]    _zz_ctrl_52;
  wire       [3:0]    _zz_ctrl_53;
  wire                _zz_ctrl_54;
  wire       [31:0]   _zz_ctrl_55;
  wire       [0:0]    _zz_ctrl_56;
  wire       [31:0]   _zz_ctrl_57;
  wire       [31:0]   _zz_ctrl_58;
  wire       [1:0]    _zz_ctrl_59;
  wire                _zz_ctrl_60;
  wire       [31:0]   _zz_ctrl_61;
  wire                _zz_ctrl_62;
  wire       [31:0]   _zz_ctrl_63;
  wire       [16:0]   _zz_ctrl_64;
  wire                _zz_ctrl_65;
  wire       [0:0]    _zz_ctrl_66;
  wire       [31:0]   _zz_ctrl_67;
  wire       [31:0]   _zz_ctrl_68;
  wire       [3:0]    _zz_ctrl_69;
  wire                _zz_ctrl_70;
  wire       [31:0]   _zz_ctrl_71;
  wire       [0:0]    _zz_ctrl_72;
  wire       [31:0]   _zz_ctrl_73;
  wire       [31:0]   _zz_ctrl_74;
  wire       [1:0]    _zz_ctrl_75;
  wire                _zz_ctrl_76;
  wire       [31:0]   _zz_ctrl_77;
  wire                _zz_ctrl_78;
  wire       [31:0]   _zz_ctrl_79;
  wire       [0:0]    _zz_ctrl_80;
  wire       [5:0]    _zz_ctrl_81;
  wire                _zz_ctrl_82;
  wire       [31:0]   _zz_ctrl_83;
  wire       [0:0]    _zz_ctrl_84;
  wire       [31:0]   _zz_ctrl_85;
  wire       [31:0]   _zz_ctrl_86;
  wire       [3:0]    _zz_ctrl_87;
  wire                _zz_ctrl_88;
  wire       [31:0]   _zz_ctrl_89;
  wire       [0:0]    _zz_ctrl_90;
  wire       [31:0]   _zz_ctrl_91;
  wire       [31:0]   _zz_ctrl_92;
  wire       [1:0]    _zz_ctrl_93;
  wire                _zz_ctrl_94;
  wire       [31:0]   _zz_ctrl_95;
  wire                _zz_ctrl_96;
  wire       [31:0]   _zz_ctrl_97;
  wire       [14:0]   _zz_ctrl_98;
  wire                _zz_ctrl_99;
  wire       [0:0]    _zz_ctrl_100;
  wire       [31:0]   _zz_ctrl_101;
  wire       [31:0]   _zz_ctrl_102;
  wire       [0:0]    _zz_ctrl_103;
  wire       [31:0]   _zz_ctrl_104;
  wire       [31:0]   _zz_ctrl_105;
  wire       [0:0]    _zz_ctrl_106;
  wire       [1:0]    _zz_ctrl_107;
  wire                _zz_ctrl_108;
  wire       [31:0]   _zz_ctrl_109;
  wire                _zz_ctrl_110;
  wire       [31:0]   _zz_ctrl_111;
  wire       [12:0]   _zz_ctrl_112;
  wire                _zz_ctrl_113;
  wire       [0:0]    _zz_ctrl_114;
  wire       [31:0]   _zz_ctrl_115;
  wire       [31:0]   _zz_ctrl_116;
  wire       [1:0]    _zz_ctrl_117;
  wire                _zz_ctrl_118;
  wire       [31:0]   _zz_ctrl_119;
  wire                _zz_ctrl_120;
  wire       [31:0]   _zz_ctrl_121;
  wire       [0:0]    _zz_ctrl_122;
  wire       [3:0]    _zz_ctrl_123;
  wire                _zz_ctrl_124;
  wire       [31:0]   _zz_ctrl_125;
  wire       [0:0]    _zz_ctrl_126;
  wire       [31:0]   _zz_ctrl_127;
  wire       [31:0]   _zz_ctrl_128;
  wire       [1:0]    _zz_ctrl_129;
  wire                _zz_ctrl_130;
  wire       [31:0]   _zz_ctrl_131;
  wire                _zz_ctrl_132;
  wire       [31:0]   _zz_ctrl_133;
  wire       [10:0]   _zz_ctrl_134;
  wire                _zz_ctrl_135;
  wire       [0:0]    _zz_ctrl_136;
  wire       [31:0]   _zz_ctrl_137;
  wire       [31:0]   _zz_ctrl_138;
  wire       [2:0]    _zz_ctrl_139;
  wire                _zz_ctrl_140;
  wire       [31:0]   _zz_ctrl_141;
  wire       [0:0]    _zz_ctrl_142;
  wire       [31:0]   _zz_ctrl_143;
  wire       [31:0]   _zz_ctrl_144;
  wire       [0:0]    _zz_ctrl_145;
  wire       [31:0]   _zz_ctrl_146;
  wire       [31:0]   _zz_ctrl_147;
  wire       [0:0]    _zz_ctrl_148;
  wire       [3:0]    _zz_ctrl_149;
  wire                _zz_ctrl_150;
  wire       [31:0]   _zz_ctrl_151;
  wire       [0:0]    _zz_ctrl_152;
  wire       [31:0]   _zz_ctrl_153;
  wire       [31:0]   _zz_ctrl_154;
  wire       [1:0]    _zz_ctrl_155;
  wire                _zz_ctrl_156;
  wire       [31:0]   _zz_ctrl_157;
  wire                _zz_ctrl_158;
  wire       [31:0]   _zz_ctrl_159;
  wire       [8:0]    _zz_ctrl_160;
  wire                _zz_ctrl_161;
  wire       [0:0]    _zz_ctrl_162;
  wire       [31:0]   _zz_ctrl_163;
  wire       [31:0]   _zz_ctrl_164;
  wire       [4:0]    _zz_ctrl_165;
  wire                _zz_ctrl_166;
  wire       [31:0]   _zz_ctrl_167;
  wire       [0:0]    _zz_ctrl_168;
  wire       [31:0]   _zz_ctrl_169;
  wire       [31:0]   _zz_ctrl_170;
  wire       [2:0]    _zz_ctrl_171;
  wire                _zz_ctrl_172;
  wire       [31:0]   _zz_ctrl_173;
  wire       [0:0]    _zz_ctrl_174;
  wire       [31:0]   _zz_ctrl_175;
  wire       [31:0]   _zz_ctrl_176;
  wire       [0:0]    _zz_ctrl_177;
  wire       [31:0]   _zz_ctrl_178;
  wire       [31:0]   _zz_ctrl_179;
  wire       [0:0]    _zz_ctrl_180;
  wire       [4:0]    _zz_ctrl_181;
  wire                _zz_ctrl_182;
  wire       [31:0]   _zz_ctrl_183;
  wire       [0:0]    _zz_ctrl_184;
  wire       [31:0]   _zz_ctrl_185;
  wire       [31:0]   _zz_ctrl_186;
  wire       [2:0]    _zz_ctrl_187;
  wire                _zz_ctrl_188;
  wire       [31:0]   _zz_ctrl_189;
  wire       [0:0]    _zz_ctrl_190;
  wire       [31:0]   _zz_ctrl_191;
  wire       [31:0]   _zz_ctrl_192;
  wire       [0:0]    _zz_ctrl_193;
  wire       [31:0]   _zz_ctrl_194;
  wire       [31:0]   _zz_ctrl_195;
  wire       [6:0]    _zz_ctrl_196;
  wire                _zz_ctrl_197;
  wire                _zz_ctrl_198;
  wire       [31:0]   _zz_ctrl_199;
  wire       [0:0]    _zz_ctrl_200;
  wire       [0:0]    _zz_ctrl_201;
  wire       [31:0]   _zz_ctrl_202;
  wire       [31:0]   _zz_ctrl_203;
  wire       [4:0]    _zz_ctrl_204;
  wire                _zz_ctrl_205;
  wire       [0:0]    _zz_ctrl_206;
  wire       [31:0]   _zz_ctrl_207;
  wire       [31:0]   _zz_ctrl_208;
  wire       [0:0]    _zz_ctrl_209;
  wire       [31:0]   _zz_ctrl_210;
  wire       [31:0]   _zz_ctrl_211;
  wire       [0:0]    _zz_ctrl_212;
  wire       [0:0]    _zz_ctrl_213;
  wire       [31:0]   _zz_ctrl_214;
  wire       [31:0]   _zz_ctrl_215;
  wire       [2:0]    _zz_ctrl_216;
  wire                _zz_ctrl_217;
  wire                _zz_ctrl_218;
  wire       [0:0]    _zz_ctrl_219;
  wire       [3:0]    _zz_ctrl_220;
  wire       [31:0]   _zz_ctrl_221;
  wire       [31:0]   _zz_ctrl_222;
  wire       [31:0]   _zz_ctrl_223;
  wire                _zz_ctrl_224;
  wire                _zz_ctrl_225;
  wire       [0:0]    _zz_ctrl_226;
  wire       [2:0]    _zz_ctrl_227;
  wire       [31:0]   _zz_ctrl_228;
  wire       [31:0]   _zz_ctrl_229;
  wire       [31:0]   _zz_ctrl_230;
  wire       [31:0]   _zz_ctrl_231;
  wire       [31:0]   _zz_ctrl_232;
  wire       [31:0]   _zz_fixInvalidInst;
  wire       [31:0]   _zz_fixInvalidInst_1;
  wire       [31:0]   _zz_fixInvalidInst_2;
  wire                _zz_fixInvalidInst_3;
  wire       [0:0]    _zz_fixInvalidInst_4;
  wire       [20:0]   _zz_fixInvalidInst_5;
  wire       [31:0]   _zz_fixInvalidInst_6;
  wire       [31:0]   _zz_fixInvalidInst_7;
  wire       [31:0]   _zz_fixInvalidInst_8;
  wire                _zz_fixInvalidInst_9;
  wire       [0:0]    _zz_fixInvalidInst_10;
  wire       [14:0]   _zz_fixInvalidInst_11;
  wire       [31:0]   _zz_fixInvalidInst_12;
  wire       [31:0]   _zz_fixInvalidInst_13;
  wire       [31:0]   _zz_fixInvalidInst_14;
  wire                _zz_fixInvalidInst_15;
  wire       [0:0]    _zz_fixInvalidInst_16;
  wire       [8:0]    _zz_fixInvalidInst_17;
  wire       [31:0]   _zz_fixInvalidInst_18;
  wire       [31:0]   _zz_fixInvalidInst_19;
  wire       [31:0]   _zz_fixInvalidInst_20;
  wire                _zz_fixInvalidInst_21;
  wire       [0:0]    _zz_fixInvalidInst_22;
  wire       [2:0]    _zz_fixInvalidInst_23;
  wire       [25:0]   ctrl;
  wire       [57:0]   fixDebug;
  wire       [58:0]   fixInvalidInst;

  assign _zz_ctrl = 32'h70000000;
  assign _zz_ctrl_1 = ((instr_i & 32'h50000000) == 32'h10000000);
  assign _zz_ctrl_2 = ((instr_i & _zz_ctrl_3) == 32'h40000000);
  assign _zz_ctrl_4 = {(_zz_ctrl_5 == _zz_ctrl_6),{_zz_ctrl_7,{_zz_ctrl_9,_zz_ctrl_12}}};
  assign _zz_ctrl_15 = ((instr_i & _zz_ctrl_16) == 32'h40000000);
  assign _zz_ctrl_17 = ((instr_i & _zz_ctrl_18) == 32'h40000000);
  assign _zz_ctrl_19 = ((instr_i & _zz_ctrl_20) == 32'h60000000);
  assign _zz_ctrl_21 = (|{_zz_ctrl_22,_zz_ctrl_24});
  assign _zz_ctrl_26 = (|_zz_ctrl_27);
  assign _zz_ctrl_29 = {(|_zz_ctrl_30),{_zz_ctrl_39,{_zz_ctrl_52,_zz_ctrl_64}}};
  assign _zz_ctrl_3 = 32'h58000000;
  assign _zz_ctrl_5 = (instr_i & 32'h66c00000);
  assign _zz_ctrl_6 = 32'h02000000;
  assign _zz_ctrl_7 = ((instr_i & _zz_ctrl_8) == 32'h00200000);
  assign _zz_ctrl_9 = (_zz_ctrl_10 == _zz_ctrl_11);
  assign _zz_ctrl_12 = (_zz_ctrl_13 == _zz_ctrl_14);
  assign _zz_ctrl_16 = 32'h70000000;
  assign _zz_ctrl_18 = 32'h68000000;
  assign _zz_ctrl_20 = 32'h60000000;
  assign _zz_ctrl_22 = ((instr_i & _zz_ctrl_23) == 32'h24000000);
  assign _zz_ctrl_24 = ((instr_i & _zz_ctrl_25) == 32'h5c000000);
  assign _zz_ctrl_27 = ((instr_i & _zz_ctrl_28) == 32'h00200000);
  assign _zz_ctrl_30 = {_zz_ctrl_31,{_zz_ctrl_33,_zz_ctrl_36}};
  assign _zz_ctrl_39 = (|{_zz_ctrl_40,_zz_ctrl_43});
  assign _zz_ctrl_52 = (|_zz_ctrl_53);
  assign _zz_ctrl_64 = {_zz_ctrl_65,{_zz_ctrl_80,_zz_ctrl_98}};
  assign _zz_ctrl_8 = 32'h66290000;
  assign _zz_ctrl_10 = (instr_i & 32'h66290000);
  assign _zz_ctrl_11 = 32'h00080000;
  assign _zz_ctrl_13 = (instr_i & 32'h66268000);
  assign _zz_ctrl_14 = 32'h00020000;
  assign _zz_ctrl_23 = 32'h24000000;
  assign _zz_ctrl_25 = 32'h5c000000;
  assign _zz_ctrl_28 = 32'h66280000;
  assign _zz_ctrl_31 = ((instr_i & _zz_ctrl_32) == 32'h00090000);
  assign _zz_ctrl_33 = (_zz_ctrl_34 == _zz_ctrl_35);
  assign _zz_ctrl_36 = (_zz_ctrl_37 == _zz_ctrl_38);
  assign _zz_ctrl_40 = (_zz_ctrl_41 == _zz_ctrl_42);
  assign _zz_ctrl_43 = {_zz_ctrl_44,{_zz_ctrl_46,_zz_ctrl_49}};
  assign _zz_ctrl_53 = {_zz_ctrl_54,{_zz_ctrl_56,_zz_ctrl_59}};
  assign _zz_ctrl_65 = (|{_zz_ctrl_66,_zz_ctrl_69});
  assign _zz_ctrl_80 = (|_zz_ctrl_81);
  assign _zz_ctrl_98 = {_zz_ctrl_99,{_zz_ctrl_106,_zz_ctrl_112}};
  assign _zz_ctrl_32 = 32'h66290000;
  assign _zz_ctrl_34 = (instr_i & 32'h66488000);
  assign _zz_ctrl_35 = 32'h00088000;
  assign _zz_ctrl_37 = (instr_i & 32'h66508000);
  assign _zz_ctrl_38 = 32'h00008000;
  assign _zz_ctrl_41 = (instr_i & 32'h58000000);
  assign _zz_ctrl_42 = 32'h10000000;
  assign _zz_ctrl_44 = ((instr_i & _zz_ctrl_45) == 32'h00040000);
  assign _zz_ctrl_46 = (_zz_ctrl_47 == _zz_ctrl_48);
  assign _zz_ctrl_49 = (_zz_ctrl_50 == _zz_ctrl_51);
  assign _zz_ctrl_54 = ((instr_i & _zz_ctrl_55) == 32'h01800000);
  assign _zz_ctrl_56 = (_zz_ctrl_57 == _zz_ctrl_58);
  assign _zz_ctrl_59 = {_zz_ctrl_60,_zz_ctrl_62};
  assign _zz_ctrl_66 = (_zz_ctrl_67 == _zz_ctrl_68);
  assign _zz_ctrl_69 = {_zz_ctrl_70,{_zz_ctrl_72,_zz_ctrl_75}};
  assign _zz_ctrl_81 = {_zz_ctrl_82,{_zz_ctrl_84,_zz_ctrl_87}};
  assign _zz_ctrl_99 = (|{_zz_ctrl_100,_zz_ctrl_103});
  assign _zz_ctrl_106 = (|_zz_ctrl_107);
  assign _zz_ctrl_112 = {_zz_ctrl_113,{_zz_ctrl_122,_zz_ctrl_134}};
  assign _zz_ctrl_45 = 32'h66140000;
  assign _zz_ctrl_47 = (instr_i & 32'h66068000);
  assign _zz_ctrl_48 = 32'h00068000;
  assign _zz_ctrl_50 = (instr_i & 32'h662c0000);
  assign _zz_ctrl_51 = 32'h00080000;
  assign _zz_ctrl_55 = 32'h71800000;
  assign _zz_ctrl_57 = (instr_i & 32'h664c0000);
  assign _zz_ctrl_58 = 32'h00400000;
  assign _zz_ctrl_60 = ((instr_i & _zz_ctrl_61) == 32'h00040000);
  assign _zz_ctrl_62 = ((instr_i & _zz_ctrl_63) == 32'h00050000);
  assign _zz_ctrl_67 = (instr_i & 32'h66800000);
  assign _zz_ctrl_68 = 32'h02000000;
  assign _zz_ctrl_70 = ((instr_i & _zz_ctrl_71) == 32'h00020000);
  assign _zz_ctrl_72 = (_zz_ctrl_73 == _zz_ctrl_74);
  assign _zz_ctrl_75 = {_zz_ctrl_76,_zz_ctrl_78};
  assign _zz_ctrl_82 = ((instr_i & _zz_ctrl_83) == 32'h10000000);
  assign _zz_ctrl_84 = (_zz_ctrl_85 == _zz_ctrl_86);
  assign _zz_ctrl_87 = {_zz_ctrl_88,{_zz_ctrl_90,_zz_ctrl_93}};
  assign _zz_ctrl_100 = (_zz_ctrl_101 == _zz_ctrl_102);
  assign _zz_ctrl_103 = (_zz_ctrl_104 == _zz_ctrl_105);
  assign _zz_ctrl_107 = {_zz_ctrl_108,_zz_ctrl_110};
  assign _zz_ctrl_113 = (|{_zz_ctrl_114,_zz_ctrl_117});
  assign _zz_ctrl_122 = (|_zz_ctrl_123);
  assign _zz_ctrl_134 = {_zz_ctrl_135,{_zz_ctrl_148,_zz_ctrl_160}};
  assign _zz_ctrl_61 = 32'h660c8000;
  assign _zz_ctrl_63 = 32'h660f0000;
  assign _zz_ctrl_71 = 32'h66260000;
  assign _zz_ctrl_73 = (instr_i & 32'h66228000);
  assign _zz_ctrl_74 = 32'h00020000;
  assign _zz_ctrl_76 = ((instr_i & _zz_ctrl_77) == 32'h00400000);
  assign _zz_ctrl_78 = ((instr_i & _zz_ctrl_79) == 32'h00040000);
  assign _zz_ctrl_83 = 32'h58000000;
  assign _zz_ctrl_85 = (instr_i & 32'h71400000);
  assign _zz_ctrl_86 = 32'h01400000;
  assign _zz_ctrl_88 = ((instr_i & _zz_ctrl_89) == 32'h00060000);
  assign _zz_ctrl_90 = (_zz_ctrl_91 == _zz_ctrl_92);
  assign _zz_ctrl_93 = {_zz_ctrl_94,_zz_ctrl_96};
  assign _zz_ctrl_101 = (instr_i & 32'h64400000);
  assign _zz_ctrl_102 = 32'h00400000;
  assign _zz_ctrl_104 = (instr_i & 32'h66000000);
  assign _zz_ctrl_105 = 32'h02000000;
  assign _zz_ctrl_108 = ((instr_i & _zz_ctrl_109) == 32'h10000000);
  assign _zz_ctrl_110 = ((instr_i & _zz_ctrl_111) == 32'h40000000);
  assign _zz_ctrl_114 = (_zz_ctrl_115 == _zz_ctrl_116);
  assign _zz_ctrl_117 = {_zz_ctrl_118,_zz_ctrl_120};
  assign _zz_ctrl_123 = {_zz_ctrl_124,{_zz_ctrl_126,_zz_ctrl_129}};
  assign _zz_ctrl_135 = (|{_zz_ctrl_136,_zz_ctrl_139});
  assign _zz_ctrl_148 = (|_zz_ctrl_149);
  assign _zz_ctrl_160 = {_zz_ctrl_161,{_zz_ctrl_180,_zz_ctrl_196}};
  assign _zz_ctrl_77 = 32'h664c0000;
  assign _zz_ctrl_79 = 32'h664d0000;
  assign _zz_ctrl_89 = 32'h66068000;
  assign _zz_ctrl_91 = (instr_i & 32'h66250000);
  assign _zz_ctrl_92 = 32'h00010000;
  assign _zz_ctrl_94 = ((instr_i & _zz_ctrl_95) == 32'h00400000);
  assign _zz_ctrl_96 = ((instr_i & _zz_ctrl_97) == 32'h00008000);
  assign _zz_ctrl_109 = 32'h10000000;
  assign _zz_ctrl_111 = 32'h40000000;
  assign _zz_ctrl_115 = (instr_i & 32'h68000000);
  assign _zz_ctrl_116 = 32'h08000000;
  assign _zz_ctrl_118 = ((instr_i & _zz_ctrl_119) == 32'h40000000);
  assign _zz_ctrl_120 = ((instr_i & _zz_ctrl_121) == 32'h02000000);
  assign _zz_ctrl_124 = ((instr_i & _zz_ctrl_125) == 32'h04000000);
  assign _zz_ctrl_126 = (_zz_ctrl_127 == _zz_ctrl_128);
  assign _zz_ctrl_129 = {_zz_ctrl_130,_zz_ctrl_132};
  assign _zz_ctrl_136 = (_zz_ctrl_137 == _zz_ctrl_138);
  assign _zz_ctrl_139 = {_zz_ctrl_140,{_zz_ctrl_142,_zz_ctrl_145}};
  assign _zz_ctrl_149 = {_zz_ctrl_150,{_zz_ctrl_152,_zz_ctrl_155}};
  assign _zz_ctrl_161 = (|{_zz_ctrl_162,_zz_ctrl_165});
  assign _zz_ctrl_180 = (|_zz_ctrl_181);
  assign _zz_ctrl_196 = {_zz_ctrl_197,{_zz_ctrl_200,_zz_ctrl_204}};
  assign _zz_ctrl_95 = 32'h664c0000;
  assign _zz_ctrl_97 = 32'h666a8000;
  assign _zz_ctrl_119 = 32'h68000000;
  assign _zz_ctrl_121 = 32'h47000000;
  assign _zz_ctrl_125 = 32'h44000000;
  assign _zz_ctrl_127 = (instr_i & 32'h41000000);
  assign _zz_ctrl_128 = 32'h01000000;
  assign _zz_ctrl_130 = ((instr_i & _zz_ctrl_131) == 32'h20000000);
  assign _zz_ctrl_132 = ((instr_i & _zz_ctrl_133) == 32'h00000000);
  assign _zz_ctrl_137 = (instr_i & 32'h46408000);
  assign _zz_ctrl_138 = 32'h06408000;
  assign _zz_ctrl_140 = ((instr_i & _zz_ctrl_141) == 32'h06401800);
  assign _zz_ctrl_142 = (_zz_ctrl_143 == _zz_ctrl_144);
  assign _zz_ctrl_145 = (_zz_ctrl_146 == _zz_ctrl_147);
  assign _zz_ctrl_150 = ((instr_i & _zz_ctrl_151) == 32'h06400000);
  assign _zz_ctrl_152 = (_zz_ctrl_153 == _zz_ctrl_154);
  assign _zz_ctrl_155 = {_zz_ctrl_156,_zz_ctrl_158};
  assign _zz_ctrl_162 = (_zz_ctrl_163 == _zz_ctrl_164);
  assign _zz_ctrl_165 = {_zz_ctrl_166,{_zz_ctrl_168,_zz_ctrl_171}};
  assign _zz_ctrl_181 = {_zz_ctrl_182,{_zz_ctrl_184,_zz_ctrl_187}};
  assign _zz_ctrl_197 = (|_zz_ctrl_198);
  assign _zz_ctrl_200 = (|_zz_ctrl_201);
  assign _zz_ctrl_204 = {_zz_ctrl_205,{_zz_ctrl_212,_zz_ctrl_216}};
  assign _zz_ctrl_131 = 32'h62000000;
  assign _zz_ctrl_133 = 32'h42400000;
  assign _zz_ctrl_141 = 32'h46401800;
  assign _zz_ctrl_143 = (instr_i & 32'h66580000);
  assign _zz_ctrl_144 = 32'h00080000;
  assign _zz_ctrl_146 = (instr_i & 32'h66700000);
  assign _zz_ctrl_147 = 32'h00000000;
  assign _zz_ctrl_151 = 32'h46408800;
  assign _zz_ctrl_153 = (instr_i & 32'h46409000);
  assign _zz_ctrl_154 = 32'h06400000;
  assign _zz_ctrl_156 = ((instr_i & _zz_ctrl_157) == 32'h00000000);
  assign _zz_ctrl_158 = ((instr_i & _zz_ctrl_159) == 32'h00080000);
  assign _zz_ctrl_163 = (instr_i & 32'h56000000);
  assign _zz_ctrl_164 = 32'h04000000;
  assign _zz_ctrl_166 = ((instr_i & _zz_ctrl_167) == 32'h04000000);
  assign _zz_ctrl_168 = (_zz_ctrl_169 == _zz_ctrl_170);
  assign _zz_ctrl_171 = {_zz_ctrl_172,{_zz_ctrl_174,_zz_ctrl_177}};
  assign _zz_ctrl_182 = ((instr_i & _zz_ctrl_183) == 32'h06000000);
  assign _zz_ctrl_184 = (_zz_ctrl_185 == _zz_ctrl_186);
  assign _zz_ctrl_187 = {_zz_ctrl_188,{_zz_ctrl_190,_zz_ctrl_193}};
  assign _zz_ctrl_198 = ((instr_i & _zz_ctrl_199) == 32'h22400000);
  assign _zz_ctrl_201 = (_zz_ctrl_202 == _zz_ctrl_203);
  assign _zz_ctrl_205 = (|{_zz_ctrl_206,_zz_ctrl_209});
  assign _zz_ctrl_212 = (|_zz_ctrl_213);
  assign _zz_ctrl_216 = {_zz_ctrl_217,{_zz_ctrl_219,_zz_ctrl_226}};
  assign _zz_ctrl_157 = 32'h66700000;
  assign _zz_ctrl_159 = 32'h66590000;
  assign _zz_ctrl_167 = 32'h54400000;
  assign _zz_ctrl_169 = (instr_i & 32'h54018000);
  assign _zz_ctrl_170 = 32'h04008000;
  assign _zz_ctrl_172 = ((instr_i & _zz_ctrl_173) == 32'h04000000);
  assign _zz_ctrl_174 = (_zz_ctrl_175 == _zz_ctrl_176);
  assign _zz_ctrl_177 = (_zz_ctrl_178 == _zz_ctrl_179);
  assign _zz_ctrl_183 = 32'h46400000;
  assign _zz_ctrl_185 = (instr_i & 32'h46008400);
  assign _zz_ctrl_186 = 32'h06000400;
  assign _zz_ctrl_188 = ((instr_i & _zz_ctrl_189) == 32'h06001800);
  assign _zz_ctrl_190 = (_zz_ctrl_191 == _zz_ctrl_192);
  assign _zz_ctrl_193 = (_zz_ctrl_194 == _zz_ctrl_195);
  assign _zz_ctrl_199 = 32'h62400000;
  assign _zz_ctrl_202 = (instr_i & 32'h00000000);
  assign _zz_ctrl_203 = 32'h00000000;
  assign _zz_ctrl_206 = (_zz_ctrl_207 == _zz_ctrl_208);
  assign _zz_ctrl_209 = (_zz_ctrl_210 == _zz_ctrl_211);
  assign _zz_ctrl_213 = (_zz_ctrl_214 == _zz_ctrl_215);
  assign _zz_ctrl_217 = (|_zz_ctrl_218);
  assign _zz_ctrl_219 = (|_zz_ctrl_220);
  assign _zz_ctrl_226 = (|_zz_ctrl_227);
  assign _zz_ctrl_173 = 32'h54010800;
  assign _zz_ctrl_175 = (instr_i & 32'h72190000);
  assign _zz_ctrl_176 = 32'h00090000;
  assign _zz_ctrl_178 = (instr_i & 32'h72700400);
  assign _zz_ctrl_179 = 32'h00000400;
  assign _zz_ctrl_189 = 32'h46009800;
  assign _zz_ctrl_191 = (instr_i & 32'h66190000);
  assign _zz_ctrl_192 = 32'h00090000;
  assign _zz_ctrl_194 = (instr_i & 32'h66700400);
  assign _zz_ctrl_195 = 32'h00000000;
  assign _zz_ctrl_207 = (instr_i & 32'h62400000);
  assign _zz_ctrl_208 = 32'h20400000;
  assign _zz_ctrl_210 = (instr_i & 32'h62400000);
  assign _zz_ctrl_211 = 32'h22000000;
  assign _zz_ctrl_214 = (instr_i & 32'h53000000);
  assign _zz_ctrl_215 = 32'h01000000;
  assign _zz_ctrl_218 = ((instr_i & 32'h60000000) == 32'h20000000);
  assign _zz_ctrl_220 = {((instr_i & _zz_ctrl_221) == 32'h40000000),{(_zz_ctrl_222 == _zz_ctrl_223),{_zz_ctrl_224,_zz_ctrl_225}}};
  assign _zz_ctrl_227 = {((instr_i & _zz_ctrl_228) == 32'h04000000),{(_zz_ctrl_229 == _zz_ctrl_230),(_zz_ctrl_231 == _zz_ctrl_232)}};
  assign _zz_ctrl_221 = 32'h40000000;
  assign _zz_ctrl_222 = (instr_i & 32'h14000000);
  assign _zz_ctrl_223 = 32'h04000000;
  assign _zz_ctrl_224 = ((instr_i & 32'h32580000) == 32'h00080000);
  assign _zz_ctrl_225 = ((instr_i & 32'h32700000) == 32'h00000000);
  assign _zz_ctrl_228 = 32'h54000000;
  assign _zz_ctrl_229 = (instr_i & 32'h720c0000);
  assign _zz_ctrl_230 = 32'h000c0000;
  assign _zz_ctrl_231 = (instr_i & 32'h72500000);
  assign _zz_ctrl_232 = 32'h00000000;
  assign _zz_fixInvalidInst = 32'hdc000000;
  assign _zz_fixInvalidInst_1 = (instr_i & 32'hf6000000);
  assign _zz_fixInvalidInst_2 = 32'h14000000;
  assign _zz_fixInvalidInst_3 = ((instr_i & 32'hfd800000) == 32'h28000000);
  assign _zz_fixInvalidInst_4 = ((instr_i & 32'hfe400000) == 32'h28000000);
  assign _zz_fixInvalidInst_5 = {((instr_i & 32'hfe800000) == 32'h28000000),{((instr_i & 32'hff000000) == 32'h04000000),{((instr_i & _zz_fixInvalidInst_6) == 32'h03400000),{(_zz_fixInvalidInst_7 == _zz_fixInvalidInst_8),{_zz_fixInvalidInst_9,{_zz_fixInvalidInst_10,_zz_fixInvalidInst_11}}}}}};
  assign _zz_fixInvalidInst_6 = 32'hff400000;
  assign _zz_fixInvalidInst_7 = (instr_i & 32'hfec00000);
  assign _zz_fixInvalidInst_8 = 32'h02800000;
  assign _zz_fixInvalidInst_9 = ((instr_i & 32'hfec00000) == 32'h02400000);
  assign _zz_fixInvalidInst_10 = ((instr_i & 32'hfbc00000) == 32'h02000000);
  assign _zz_fixInvalidInst_11 = {((instr_i & 32'hfffd0000) == 32'h00150000),{((instr_i & 32'hfff68000) == 32'h00140000),{((instr_i & _zz_fixInvalidInst_12) == 32'h00140000),{(_zz_fixInvalidInst_13 == _zz_fixInvalidInst_14),{_zz_fixInvalidInst_15,{_zz_fixInvalidInst_16,_zz_fixInvalidInst_17}}}}}};
  assign _zz_fixInvalidInst_12 = 32'hfff70000;
  assign _zz_fixInvalidInst_13 = (instr_i & 32'hfffe0000);
  assign _zz_fixInvalidInst_14 = 32'h00200000;
  assign _zz_fixInvalidInst_15 = ((instr_i & 32'hfff38000) == 32'h00100000);
  assign _zz_fixInvalidInst_16 = ((instr_i & 32'hfffa8000) == 32'h00100000);
  assign _zz_fixInvalidInst_17 = {((instr_i & 32'hfffe8000) == 32'h06488000),{((instr_i & 32'hfffe8000) == 32'h002a0000),{((instr_i & _zz_fixInvalidInst_18) == 32'h00408000),{(_zz_fixInvalidInst_19 == _zz_fixInvalidInst_20),{_zz_fixInvalidInst_21,{_zz_fixInvalidInst_22,_zz_fixInvalidInst_23}}}}}};
  assign _zz_fixInvalidInst_18 = 32'hfffb8000;
  assign _zz_fixInvalidInst_19 = (instr_i & 32'hfff78000);
  assign _zz_fixInvalidInst_20 = 32'h00408000;
  assign _zz_fixInvalidInst_21 = ((instr_i & 32'hffff0000) == 32'h00120000);
  assign _zz_fixInvalidInst_22 = ((instr_i & 32'hfffff800) == 32'h06483000);
  assign _zz_fixInvalidInst_23 = {((instr_i & 32'hfffff400) == 32'h06483000),{((instr_i & 32'hfffff800) == 32'h06482800),((instr_i & 32'hfffff800) == 32'h00006000)}};
  assign ctrl = {(|((instr_i & _zz_ctrl) == 32'h40000000)),{(|{_zz_ctrl_1,{_zz_ctrl_2,_zz_ctrl_4}}),{(|{_zz_ctrl_15,_zz_ctrl_17}),{(|_zz_ctrl_19),{_zz_ctrl_21,{_zz_ctrl_26,_zz_ctrl_29}}}}}};
  assign fixDebug = {instr_i,ctrl};
  assign fixInvalidInst = {fixDebug,(! (|{((instr_i & 32'hf0000000) == 32'h50000000),{((instr_i & 32'hf0000000) == 32'h60000000),{((instr_i & _zz_fixInvalidInst) == 32'h4c000000),{(_zz_fixInvalidInst_1 == _zz_fixInvalidInst_2),{_zz_fixInvalidInst_3,{_zz_fixInvalidInst_4,_zz_fixInvalidInst_5}}}}}}))};
  assign option_code_o = fixInvalidInst;

endmodule


