// ==============================================================================
// Copyright (c) 2014-2024 All rights reserved
// ==============================================================================
// Author  : SuYang 2506806016@qq.com
// File    : Level2TranslationLookasideBuffer.sv
// Create  : 2024-03-01 22:21:08
// Revise  : 2024-03-01 22:21:08
// Description :
//   L2 TLB
// Parameter   :
//   ...
//   ...
// IO Port     :
//   ...
//   ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
// -----------------------------------------------------------------------------
// xx-xx-xx |            |     0.1     |    Original Version
// ...
// ==============================================================================

module Level2TranslationLookasideBuffer (
  input clk,    // Clock
  input rst_n,  // Asynchronous reset active low
  
);

endmodule : Level2TranslationLookasideBuffer

